module And(
  input a,b,c,d,
  output s);
  
  assign s = a&b&c&d;
  
endmodule