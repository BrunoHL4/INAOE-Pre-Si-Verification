module Not_Gate(
   input a,
  output c);
  
  assign c = ~a;
  
endmodule