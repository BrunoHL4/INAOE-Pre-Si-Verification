module And_3(
   input a,b,c,
  output s);
  
  assign s = a&b&c;
  
endmodule