module SegmentoF(a,b,c,x);
   input a,b,c;
  output x;
  
  assign x=1;
  
endmodule