module And_Gate4(
   input a,b,c,d,
  output e);
  
  assign e = a&b&c&d;
  
endmodule