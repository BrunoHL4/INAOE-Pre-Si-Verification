module And_Gate2(
   input a,b,
  output c);
  
  assign c = a&b;
  
endmodule