module Or(
   input a,b,c,
  output s);
  
  assign s = a|b|c;
  
endmodule