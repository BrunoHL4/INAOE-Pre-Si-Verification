module SegmentoD(a,b,c,x);
   input a,b,c;
  output x;
  
  assign x=~c;
  
endmodule