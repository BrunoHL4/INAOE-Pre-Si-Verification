module And_Gate3(
   input a,b,c,
  output d);
  
  assign d = a&b&c;
  
endmodule