module And_Gate(
   input a,b,
  output c);
  
  assign c = a&b;
  
endmodule