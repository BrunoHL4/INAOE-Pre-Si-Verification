module Not(
   input a,
  output s);
  
  assign s = ~a;
  
endmodule