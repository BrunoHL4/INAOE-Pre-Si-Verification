module Not(
   input a,
  output c);
  
  assign c = ~a;
  
endmodule