module Xor_Gate(
   input a,b,
  output c);
  
  assign c = a^b;
  
endmodule