module SegmentoI(a,b,c,x);
   input a,b,c;
  output x;
  
  assign x=0;
  
endmodule